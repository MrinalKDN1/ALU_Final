interface alu16_if;
 logic [15:0] a;
 logic [15:0] b;
 logic [2:0] op;
 logic [15:0] y;
  
endinterface
