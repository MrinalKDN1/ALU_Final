`include"alu_transection.sv"
`include"alu_generator.sv"
`include"alu_driver.sv"
`include"alu_monitor.sv"
`include"alu_agent.sv"
`include"alu_scoreboard.sv"
`include"alu_env.sv"
